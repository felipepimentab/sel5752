library work;
use work.riscv_pkg.all;

entity datapath is
	generic(
		Width : natural := 32
	);
	port(clk, reset: in BIT;
		ResultSrc: in BIT_VECTOR(1 downto 0);
		PCSrc, ALUSrc: in BIT;
		RegWrite: in BIT;
		ImmSrc: in BIT_VECTOR(1 downto 0);
		ALUControl: in BIT_VECTOR(2 downto 0);
		Zero: out BIT;
		PC: buffer BIT_VECTOR(Width-1 downto 0);
		Instr: in BIT_VECTOR(Width-1 downto 0);
		ALUResult, WriteData: buffer BIT_VECTOR(Width-1 downto 0);
		ReadData: in BIT_VECTOR(Width-1 downto 0));
end;

architecture struct of datapath is
	component flopr generic(width: integer);
		port(clk, reset: in BIT;
				d: in BIT_VECTOR(width-1 downto 0);
				q: out BIT_VECTOR(width-1 downto 0));
	end component;
	component adder
		port(a, b: in BIT_VECTOR(Width-1 downto 0);
				y: out BIT_VECTOR(Width-1 downto 0));
	end component;
	component mux2 generic(width: integer);
		port(d0, d1: in BIT_VECTOR(width-1 downto 0);
				s: in BIT;
				y: out BIT_VECTOR(width-1 downto 0));
	end component;
	component mux3 generic(width: integer);
		port(d0, d1, d2: in BIT_VECTOR(width-1 downto 0);
				s: in BIT_VECTOR(1 downto 0);
				y: out BIT_VECTOR(width-1 downto 0));
	end component;
	component regfile
		port(clk: in BIT;
				we3: in BIT;
				a1, a2, a3: in BIT_VECTOR(4 downto 0);
				wd3: in BIT_VECTOR(Width-1 downto 0);
				rd1, rd2: out BIT_VECTOR(Width-1 downto 0));
	end component;
	component extend
		port(instr: in BIT_VECTOR(Width-1 downto 7);
				immsrc: in BIT_VECTOR(1 downto 0);
				immext: out BIT_VECTOR(Width-1 downto 0));
	end component;
	component alu
		port(a, b: in BIT_VECTOR(Width-1 downto 0);
				ALUControl: in BIT_VECTOR(2 downto 0);
				ALUResult: buffer BIT_VECTOR(Width-1 downto 0);
				Zero: out BIT);
	end component;
	
	signal PCNext, PCPlus4, PCTarget: BIT_VECTOR(Width-1 downto 0);
	signal ImmExt: BIT_VECTOR(Width-1 downto 0);
	signal SrcA, SrcB: BIT_VECTOR(Width-1 downto 0);
	signal Result: BIT_VECTOR(Width-1 downto 0);
begin
	-- next PC logic
	pcreg: flopr generic map(Width) port map(clk, reset, PCNext, PC);
	pcadd4: adder port map(PC, X"00000004", PCPlus4);
	pcaddbranch: adder port map(PC, ImmExt, PCTarget);
	pcmux: mux2 generic map(Width) port map(PCPlus4, PCTarget, PCSrc,
											PCNext);
	-- register file logic
	rf: regfile port map(clk, RegWrite, Instr(19 downto 15),
	Instr(24 downto 20), Instr(11 downto 7),
								Result, SrcA, WriteData);
	ext: extend port map(Instr(Width-1 downto 7), ImmSrc, ImmExt);
	-- ALU logic
	srcbmux: mux2 generic map(Width) port map(WriteData, ImmExt,
											ALUSrc, SrcB);
	mainalu: alu port map(SrcA, SrcB, ALUControl, ALUResult, Zero);
	resultmux: mux3 generic map(Width) port map(ALUResult, ReadData,
												PCPlus4, ResultSrc,
												Result);
end;