---------------------------------
-- Título: aludec
-- Descrição: ALU Decoder
-- Autor: Felipe Pimenta Bernardo
-- Data: 27/06/2024
---------------------------------

entity aludec is
    port (
        
    );
end aludec;

architecture behaviour of aludec is
    begin

    end;